module angle_to_bcd_tb;



endmodule