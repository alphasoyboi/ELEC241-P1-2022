module servo_controller_unit (output logic [11:0] angle, input logic clk, input logic n_reset, input logic [31:0] input_register);



endmodule