module IC_tb;

endmodule